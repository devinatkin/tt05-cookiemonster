`timescale 1ns / 1ps

module crumb(
input wire clk,         // Clock signal
input wire rst_n,       // Active-low reset signal
input wire en,          // Enable signal
input wire rbit,        // Random bit in 1
input wire rbit2,       // Random bit in 2
output reg clk_o,       // Clock output
output reg rst_no,      // Reset output
output reg en_o,        // Enable output
output reg rbit_o       // Random bit output

);

//Internal Registers
reg [15:0] rand_num;
reg [3:0] clk_cnt;
always@(posedge clk) begin
    if (!rst_n) begin           // Reset Event
        clk_o <= 1'b0;          // Reset clock
        rst_no <= 1'b0;         // Reset reset
        rbit_o <= 1'b0;         // Reset random bit
        en_o <= 1'b0;           // Reset enable

        rand_num <= 16'h0000;      // Reset random number
        clk_cnt <= 4'h0;        // Reset clock counter
    end else if (en) begin
        clk_o <= ~clk_o;
        rst_no <= ~rst_no;
        rbit_o <= rbit ^ rbit2;
        en_o <= en;

        //Shift in new random bit
        rand_num <= {rand_num[14:0], rbit_o};

        if (clk_cnt == 4'hF) begin
            $display("Random Number: %h", rand_num);
            clk_cnt <= 4'h0;
        end else begin
            clk_cnt <= clk_cnt + 1'b1;
        end
    end
end

endmodule

// Each crumb is part of a cookie which comprises of 16 crumbs arranged in a 4x4 grid.
// Each crumb is connected to its neighbors via 2 input 'random' bits and 1 output 'random' bit.
// While random data is typically in the rbit stream it is not guaranteed to be random, and may be set to be messages.
// The LSFR is a 64 bit LSFR with a polynomial of x^64 + x^4 + x^3 + x + 1.

// I need to guarantee that valid messages are not generated by the LSFR.
